//////////////////////////////////////////////////////////////////////
// File Name:		sh_reg.vh										//
// Function:		shify register header							//
// Discribution:													//
// Auther:			Kerwin Simth									//
// Date:			2019.12.26										//
//////////////////////////////////////////////////////////////////////

`ifndef __SH_REG_HEADER__
	`define __SH_REG_HEADER__

	`define REG_WIDTH		[13:0]
	`define INIT			14'b0

`endif
