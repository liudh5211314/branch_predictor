//////////////////////////////////////////////////////////////////////
// File Name:		mux.v											//
// Function:		multiplexer										//
// Discribution:													//
// Auther:			Kerwin Simth									//
// Date:			2019.12.28										//
//////////////////////////////////////////////////////////////////////
`timescale 1ns/100ps

module mux #(parameter WIDTH = 32) (	input	[WIDTH-1:0]		d0,d1,
										input					s,
										output	[WIDTH-1:0]		y);

	assign y = s ? d1:d0;

endmodule
