//////////////////////////////////////////////////////////////////////
// File Name:		pre_set_tab.v									//
// Function:		pre_set pattern history table header			//
// Discribution:													//
// Auther:			Kerwin Simth									//
// Date:			2019.12.29										//
//////////////////////////////////////////////////////////////////////

