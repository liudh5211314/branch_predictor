//////////////////////////////////////////////////////////////////////
// File Name:		bra_his_tab.v									//
// Function:		branch history table header						//
// Discribution:													//
// Auther:			Kerwin Simth									//
// Date:			2019.12.29										//
//////////////////////////////////////////////////////////////////////

`ifndef	__BRA_TAB_HEADER__
	`define __BRA_TAB_HEADER__

	`define ADDR_WIDTH	[9:0]
	`define	DATA_WIDTH	[9:0]
	`define	DATA_DEEPTH	[1023:0]
	`define	LOOP_CONT	1024
	`define	INIT		10'b0

`endif
