//////////////////////////////////////////////////////////////////////
// File Name:		cache_tag.vh									//
// Function:		cache tag header								//
// Discribution:													//
// Auther:			Kerwin Simth									//
// Date:			2020.01.09										//
//////////////////////////////////////////////////////////////////////
`ifndef __CACHE_TAG_HEADER__

`endif
