//////////////////////////////////////////////////////////////////////
// File Name:		fin_sta_mac.vh									//
// Function:		finite state machine header						//
// Discribution:													//
// Auther:			Kerwin Simth									//
// Date:			2019.12.27										//
//////////////////////////////////////////////////////////////////////


