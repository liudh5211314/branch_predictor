//////////////////////////////////////////////////////////////////////
// File Name:		pat_tab.vh										//
// Function:		pattern history table header					//
// Discribution:													//
// Auther:			Kerwin Simth									//
// Date:			2019.12.27										//
//////////////////////////////////////////////////////////////////////

`ifndef __PAT_TAB_HEADER__
	`define __PAT_TAB_HEADER__

	`define DATA_WIDTH		[1:0]
	`define WR_ADDR			[13:0]
	`define DATA_DEEPTH		[16383:0]
	`define LOOP_TIMES		16384

	`define INIT			2'b10

`endif
