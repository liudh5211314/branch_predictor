//////////////////////////////////////////////////////////////////////
// File Name:		sel_tab.vh										//
// Function:		beanch predictor selection table header			//
// Discribution:													//
// Auther:			Kerwin Simth									//
// Date:			2019.12.29										//
//////////////////////////////////////////////////////////////////////

`ifndef __SEL_TAB_HEADER__
	`define	__SEL_TAB_HEADER__

	`define TAB_WIDTH		[1:0]
	`define TAB_ADDR		[9:0]
	`define	TAB_DEEPTH		[1023:0]
	`define	LOOP_TIMES		1024
	`define	INIT			2'b10

`endif
