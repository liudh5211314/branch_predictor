//////////////////////////////////////////////////////////////////////
// File Name:		cache_ram.vh									//
// Function:		cache ram header								//
// Discribution:													//
// Auther:			Kerwin Simth									//
// Date:			2020.01.11										//
//////////////////////////////////////////////////////////////////////
`ifndef __CACHE_RAM_HEADER__
	`define __CACHE_RAM_HEADER__

	`define ADDR_WIDTH		[9:0]
	`define DATA_WIDTH		[31:0]
	`define	DATA_DEEPTH		[1023:0]
`endif

