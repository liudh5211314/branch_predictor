//////////////////////////////////////////////////////////////////////
// File Name:		predictor_top.vh								//
// Function:		predictor top header							//
// Discribution:													//
// Auther:			Kerwin Simth									//
// Date:			2019.12.31										//
//////////////////////////////////////////////////////////////////////
